`timescale 1ns/100ps

module FreeList #(
    parameter PRF_SIZE = 64,                // ����Ĵ�������
    parameter FL_SIZE = 32,                 // Free List ��С
    parameter WIDTH = 2,                    // ÿ������෢�����ָ��
    parameter ROB_SIZE = 32                 // ���� rollback head
)(
    input  logic clock,
    input  logic reset,

    // �� Dispatch �׶����������ź�
    input  logic [WIDTH-1:0] dispatch_en,    // �Ƿ���������Ĵ���
    output logic [WIDTH-1:0][$clog2(PRF_SIZE)-1:0] free_phys_regs, // �����ȥ��PRF���

    // �� ROB (retire) ���� T_old
    input  logic [WIDTH-1:0] retire_en,
    input  logic [WIDTH-1:0][$clog2(PRF_SIZE)-1:0] retired_tags,

    // �ع�֧��
    input  logic rollback_en,
    input  logic [$clog2(FL_SIZE)-1:0] recover_head
);

    // ========================
    // ���ݽṹ
    // ========================
    logic [$clog2(PRF_SIZE)-1:0] freelist[FL_SIZE-1:0];
    logic [$clog2(FL_SIZE)-1:0] head, tail;
    logic [$clog2(FL_SIZE)-1:0] next_head, next_tail;
    logic [$clog2(PRF_SIZE)-1:0] temp_list[FL_SIZE-1:0];

    // ========================
    // ����׶Σ��� freelist ����������Ĵ���
    // ========================
    always_comb begin
        next_head = head;
        for (int i = 0; i < WIDTH; i++) begin
            if (dispatch_en[i]) begin
                free_phys_regs[i] = freelist[next_head];
                next_head = (next_head + 1) % FL_SIZE;
            end else begin
                free_phys_regs[i] = '0;
            end
        end
    end

    // ========================
    // �ύ�׶Σ��� ROB ���� T_old
    // ========================
    always_comb begin
        next_tail = tail;
        temp_list = freelist;
        for (int i = 0; i < WIDTH; i++) begin
            if (retire_en[i]) begin
                temp_list[next_tail] = retired_tags[i];
                next_tail = (next_tail + 1) % FL_SIZE;
            end
        end
    end

    // ========================
    // ʱ������߼�
    // ========================
    always_ff @(posedge clock or posedge reset) begin
        if (reset) begin
            // ��ʼ�� freelist
            for (int i = 0; i < FL_SIZE; i++) begin
                freelist[i] <= i + FL_SIZE; // ����ǰ�沿�ֱ����� ARF
            end
            head <= 0;
            tail <= 0;
        end else if (rollback_en) begin
            // �ع�ʱ�ָ�����ָ��
            head <= recover_head;
        end else begin
            head <= next_head;
            tail <= next_tail;
            freelist <= temp_list;
        end
    end

endmodule
